module detector(
input [1:0] a,b,
output eq
);
assign eq=(a==b);
endmodule